/*-
 * Copyright (c) 2018 Alexandre Joannou
 * All rights reserved.
 *
 * This software was developed by SRI International and the University of
 * Cambridge Computer Laboratory (Department of Computer Science and
 * Technology) under DARPA contract HR0011-18-C-0016 ("ECATS"), as part of the
 * DARPA SSITH research programme.
 *
 * @BERI_LICENSE_HEADER_START@
 *
 * Licensed to BERI Open Systems C.I.C. (BERI) under one or more contributor
 * license agreements.  See the NOTICE file distributed with this work for
 * additional information regarding copyright ownership.  BERI licenses this
 * file to you under the BERI Hardware-Software License, Version 1.0 (the
 * "License"); you may not use this file except in compliance with the
 * License.  You may obtain a copy of the License at:
 *
 *   http://www.beri-open-systems.org/legal/license-1-0.txt
 *
 * Unless required by applicable law or agreed to in writing, Work distributed
 * under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied.  See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * @BERI_LICENSE_HEADER_END@
 */

package AXI;

import AXI4_Common_Types :: *;
import AXI4_Types :: *;
import AXI4_AW_Utils :: *;
import AXI4_W_Utils :: *;
import AXI4_B_Utils :: *;
import AXI4_AR_Utils :: *;
import AXI4_R_Utils :: *;
import AXI4_Utils :: *;
import AXI4_Interconnect :: *;
import AXI4Lite_Types :: *;
import AXI4Lite_AW_Utils :: *;
import AXI4Lite_W_Utils :: *;
import AXI4Lite_B_Utils :: *;
import AXI4Lite_AR_Utils :: *;
import AXI4Lite_R_Utils :: *;
import AXI4Lite_Utils :: *;
import AXI4Lite_Interconnect :: *;
import AXI4_AXI4Lite_Bridges :: *;

export AXI4_Common_Types :: *;
export AXI4_Types :: *;
export AXI4_AW_Utils :: *;
export AXI4_W_Utils :: *;
export AXI4_B_Utils :: *;
export AXI4_AR_Utils :: *;
export AXI4_R_Utils :: *;
export AXI4_Utils :: *;
export AXI4_Interconnect :: *;
export AXI4Lite_Types :: *;
export AXI4Lite_AW_Utils :: *;
export AXI4Lite_W_Utils :: *;
export AXI4Lite_B_Utils :: *;
export AXI4Lite_AR_Utils :: *;
export AXI4Lite_R_Utils :: *;
export AXI4Lite_Utils :: *;
export AXI4Lite_Interconnect :: *;
export AXI4_AXI4Lite_Bridges :: *;

endpackage
